
package Types;

// 基本的な定数や型の定義
import BasicTypes::*;

// ここより下に，各人の定義を追加してください

endpackage
