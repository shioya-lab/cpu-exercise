
package Types;

// データ幅は16bit
parameter DATA_WIDTH = 16;

// データパス
typedef logic [DATA_WIDTH-1:0] DataPath;

endpackage

