//
// 減算器の検証用モジュール
//



// 基本的な型を定義したファイルの読み込み
import Types::*;


//
// 減算器の検証用のモジュール
//
module SubSim;

endmodule


